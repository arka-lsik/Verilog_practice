//4x1 mux code fo behavriol design
module mux_4x1_bh(y,S,I);
  input [3:0]I;
  input [1:0]S;
  output reg y;

  always@(*)
    case(S)
      2'b00: y=I[0];
      2'b01: y=I[1];
      2'b10: y=I[2];
      2'b11: y=I[3];
      default: $display("error");
    endcase
endmodule
